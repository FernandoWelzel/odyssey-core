//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.03 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Fri Oct 11 11:58:20 2024

module Gowin_RAM16S (dout, wre, ad, di, clk);

output [255:0] dout;
input wre;
input [4:0] ad;
input [255:0] di;
input clk;

wire ad4_inv;
wire lut_f_0;
wire lut_f_1;
wire [3:0] ram16s_inst_0_dout;
wire [7:4] ram16s_inst_1_dout;
wire [11:8] ram16s_inst_2_dout;
wire [15:12] ram16s_inst_3_dout;
wire [19:16] ram16s_inst_4_dout;
wire [23:20] ram16s_inst_5_dout;
wire [27:24] ram16s_inst_6_dout;
wire [31:28] ram16s_inst_7_dout;
wire [35:32] ram16s_inst_8_dout;
wire [39:36] ram16s_inst_9_dout;
wire [43:40] ram16s_inst_10_dout;
wire [47:44] ram16s_inst_11_dout;
wire [51:48] ram16s_inst_12_dout;
wire [55:52] ram16s_inst_13_dout;
wire [59:56] ram16s_inst_14_dout;
wire [63:60] ram16s_inst_15_dout;
wire [67:64] ram16s_inst_16_dout;
wire [71:68] ram16s_inst_17_dout;
wire [75:72] ram16s_inst_18_dout;
wire [79:76] ram16s_inst_19_dout;
wire [83:80] ram16s_inst_20_dout;
wire [87:84] ram16s_inst_21_dout;
wire [91:88] ram16s_inst_22_dout;
wire [95:92] ram16s_inst_23_dout;
wire [99:96] ram16s_inst_24_dout;
wire [103:100] ram16s_inst_25_dout;
wire [107:104] ram16s_inst_26_dout;
wire [111:108] ram16s_inst_27_dout;
wire [115:112] ram16s_inst_28_dout;
wire [119:116] ram16s_inst_29_dout;
wire [123:120] ram16s_inst_30_dout;
wire [127:124] ram16s_inst_31_dout;
wire [131:128] ram16s_inst_32_dout;
wire [135:132] ram16s_inst_33_dout;
wire [139:136] ram16s_inst_34_dout;
wire [143:140] ram16s_inst_35_dout;
wire [147:144] ram16s_inst_36_dout;
wire [151:148] ram16s_inst_37_dout;
wire [155:152] ram16s_inst_38_dout;
wire [159:156] ram16s_inst_39_dout;
wire [163:160] ram16s_inst_40_dout;
wire [167:164] ram16s_inst_41_dout;
wire [171:168] ram16s_inst_42_dout;
wire [175:172] ram16s_inst_43_dout;
wire [179:176] ram16s_inst_44_dout;
wire [183:180] ram16s_inst_45_dout;
wire [187:184] ram16s_inst_46_dout;
wire [191:188] ram16s_inst_47_dout;
wire [195:192] ram16s_inst_48_dout;
wire [199:196] ram16s_inst_49_dout;
wire [203:200] ram16s_inst_50_dout;
wire [207:204] ram16s_inst_51_dout;
wire [211:208] ram16s_inst_52_dout;
wire [215:212] ram16s_inst_53_dout;
wire [219:216] ram16s_inst_54_dout;
wire [223:220] ram16s_inst_55_dout;
wire [227:224] ram16s_inst_56_dout;
wire [231:228] ram16s_inst_57_dout;
wire [235:232] ram16s_inst_58_dout;
wire [239:236] ram16s_inst_59_dout;
wire [243:240] ram16s_inst_60_dout;
wire [247:244] ram16s_inst_61_dout;
wire [251:248] ram16s_inst_62_dout;
wire [255:252] ram16s_inst_63_dout;
wire [3:0] ram16s_inst_64_dout;
wire [7:4] ram16s_inst_65_dout;
wire [11:8] ram16s_inst_66_dout;
wire [15:12] ram16s_inst_67_dout;
wire [19:16] ram16s_inst_68_dout;
wire [23:20] ram16s_inst_69_dout;
wire [27:24] ram16s_inst_70_dout;
wire [31:28] ram16s_inst_71_dout;
wire [35:32] ram16s_inst_72_dout;
wire [39:36] ram16s_inst_73_dout;
wire [43:40] ram16s_inst_74_dout;
wire [47:44] ram16s_inst_75_dout;
wire [51:48] ram16s_inst_76_dout;
wire [55:52] ram16s_inst_77_dout;
wire [59:56] ram16s_inst_78_dout;
wire [63:60] ram16s_inst_79_dout;
wire [67:64] ram16s_inst_80_dout;
wire [71:68] ram16s_inst_81_dout;
wire [75:72] ram16s_inst_82_dout;
wire [79:76] ram16s_inst_83_dout;
wire [83:80] ram16s_inst_84_dout;
wire [87:84] ram16s_inst_85_dout;
wire [91:88] ram16s_inst_86_dout;
wire [95:92] ram16s_inst_87_dout;
wire [99:96] ram16s_inst_88_dout;
wire [103:100] ram16s_inst_89_dout;
wire [107:104] ram16s_inst_90_dout;
wire [111:108] ram16s_inst_91_dout;
wire [115:112] ram16s_inst_92_dout;
wire [119:116] ram16s_inst_93_dout;
wire [123:120] ram16s_inst_94_dout;
wire [127:124] ram16s_inst_95_dout;
wire [131:128] ram16s_inst_96_dout;
wire [135:132] ram16s_inst_97_dout;
wire [139:136] ram16s_inst_98_dout;
wire [143:140] ram16s_inst_99_dout;
wire [147:144] ram16s_inst_100_dout;
wire [151:148] ram16s_inst_101_dout;
wire [155:152] ram16s_inst_102_dout;
wire [159:156] ram16s_inst_103_dout;
wire [163:160] ram16s_inst_104_dout;
wire [167:164] ram16s_inst_105_dout;
wire [171:168] ram16s_inst_106_dout;
wire [175:172] ram16s_inst_107_dout;
wire [179:176] ram16s_inst_108_dout;
wire [183:180] ram16s_inst_109_dout;
wire [187:184] ram16s_inst_110_dout;
wire [191:188] ram16s_inst_111_dout;
wire [195:192] ram16s_inst_112_dout;
wire [199:196] ram16s_inst_113_dout;
wire [203:200] ram16s_inst_114_dout;
wire [207:204] ram16s_inst_115_dout;
wire [211:208] ram16s_inst_116_dout;
wire [215:212] ram16s_inst_117_dout;
wire [219:216] ram16s_inst_118_dout;
wire [223:220] ram16s_inst_119_dout;
wire [227:224] ram16s_inst_120_dout;
wire [231:228] ram16s_inst_121_dout;
wire [235:232] ram16s_inst_122_dout;
wire [239:236] ram16s_inst_123_dout;
wire [243:240] ram16s_inst_124_dout;
wire [247:244] ram16s_inst_125_dout;
wire [251:248] ram16s_inst_126_dout;
wire [255:252] ram16s_inst_127_dout;
wire gw_vcc;

assign gw_vcc = 1'b1;

INV inv_inst_0 (.I(ad[4]), .O(ad4_inv));

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(wre),
  .I1(ad4_inv),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_0.INIT = 16'h8000;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(wre),
  .I1(ad[4]),
  .I2(gw_vcc),
  .I3(gw_vcc)
);
defparam lut_inst_1.INIT = 16'h8000;
RAM16S4 ram16s_inst_0 (
    .DO(ram16s_inst_0_dout[3:0]),
    .DI(di[3:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_0.INIT_0 = 16'h0000;
defparam ram16s_inst_0.INIT_1 = 16'h0000;
defparam ram16s_inst_0.INIT_2 = 16'h0000;
defparam ram16s_inst_0.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_1 (
    .DO(ram16s_inst_1_dout[7:4]),
    .DI(di[7:4]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_1.INIT_0 = 16'h0000;
defparam ram16s_inst_1.INIT_1 = 16'h0000;
defparam ram16s_inst_1.INIT_2 = 16'h0000;
defparam ram16s_inst_1.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_2 (
    .DO(ram16s_inst_2_dout[11:8]),
    .DI(di[11:8]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_2.INIT_0 = 16'h0000;
defparam ram16s_inst_2.INIT_1 = 16'h0000;
defparam ram16s_inst_2.INIT_2 = 16'h0000;
defparam ram16s_inst_2.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_3 (
    .DO(ram16s_inst_3_dout[15:12]),
    .DI(di[15:12]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_3.INIT_0 = 16'h0000;
defparam ram16s_inst_3.INIT_1 = 16'h0000;
defparam ram16s_inst_3.INIT_2 = 16'h0000;
defparam ram16s_inst_3.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_4 (
    .DO(ram16s_inst_4_dout[19:16]),
    .DI(di[19:16]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_4.INIT_0 = 16'h0000;
defparam ram16s_inst_4.INIT_1 = 16'h0000;
defparam ram16s_inst_4.INIT_2 = 16'h0000;
defparam ram16s_inst_4.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_5 (
    .DO(ram16s_inst_5_dout[23:20]),
    .DI(di[23:20]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_5.INIT_0 = 16'h0000;
defparam ram16s_inst_5.INIT_1 = 16'h0000;
defparam ram16s_inst_5.INIT_2 = 16'h0000;
defparam ram16s_inst_5.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_6 (
    .DO(ram16s_inst_6_dout[27:24]),
    .DI(di[27:24]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_6.INIT_0 = 16'h0000;
defparam ram16s_inst_6.INIT_1 = 16'h0000;
defparam ram16s_inst_6.INIT_2 = 16'h0000;
defparam ram16s_inst_6.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_7 (
    .DO(ram16s_inst_7_dout[31:28]),
    .DI(di[31:28]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_7.INIT_0 = 16'h0000;
defparam ram16s_inst_7.INIT_1 = 16'h0000;
defparam ram16s_inst_7.INIT_2 = 16'h0000;
defparam ram16s_inst_7.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_8 (
    .DO(ram16s_inst_8_dout[35:32]),
    .DI(di[35:32]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_8.INIT_0 = 16'h0000;
defparam ram16s_inst_8.INIT_1 = 16'h0000;
defparam ram16s_inst_8.INIT_2 = 16'h0000;
defparam ram16s_inst_8.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_9 (
    .DO(ram16s_inst_9_dout[39:36]),
    .DI(di[39:36]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_9.INIT_0 = 16'h0000;
defparam ram16s_inst_9.INIT_1 = 16'h0000;
defparam ram16s_inst_9.INIT_2 = 16'h0000;
defparam ram16s_inst_9.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_10 (
    .DO(ram16s_inst_10_dout[43:40]),
    .DI(di[43:40]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_10.INIT_0 = 16'h0000;
defparam ram16s_inst_10.INIT_1 = 16'h0000;
defparam ram16s_inst_10.INIT_2 = 16'h0000;
defparam ram16s_inst_10.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_11 (
    .DO(ram16s_inst_11_dout[47:44]),
    .DI(di[47:44]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_11.INIT_0 = 16'h0000;
defparam ram16s_inst_11.INIT_1 = 16'h0000;
defparam ram16s_inst_11.INIT_2 = 16'h0000;
defparam ram16s_inst_11.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_12 (
    .DO(ram16s_inst_12_dout[51:48]),
    .DI(di[51:48]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_12.INIT_0 = 16'h0000;
defparam ram16s_inst_12.INIT_1 = 16'h0000;
defparam ram16s_inst_12.INIT_2 = 16'h0000;
defparam ram16s_inst_12.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_13 (
    .DO(ram16s_inst_13_dout[55:52]),
    .DI(di[55:52]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_13.INIT_0 = 16'h0000;
defparam ram16s_inst_13.INIT_1 = 16'h0000;
defparam ram16s_inst_13.INIT_2 = 16'h0000;
defparam ram16s_inst_13.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_14 (
    .DO(ram16s_inst_14_dout[59:56]),
    .DI(di[59:56]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_14.INIT_0 = 16'h0000;
defparam ram16s_inst_14.INIT_1 = 16'h0000;
defparam ram16s_inst_14.INIT_2 = 16'h0000;
defparam ram16s_inst_14.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_15 (
    .DO(ram16s_inst_15_dout[63:60]),
    .DI(di[63:60]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_15.INIT_0 = 16'h0000;
defparam ram16s_inst_15.INIT_1 = 16'h0000;
defparam ram16s_inst_15.INIT_2 = 16'h0000;
defparam ram16s_inst_15.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_16 (
    .DO(ram16s_inst_16_dout[67:64]),
    .DI(di[67:64]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_16.INIT_0 = 16'h0000;
defparam ram16s_inst_16.INIT_1 = 16'h0000;
defparam ram16s_inst_16.INIT_2 = 16'h0000;
defparam ram16s_inst_16.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_17 (
    .DO(ram16s_inst_17_dout[71:68]),
    .DI(di[71:68]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_17.INIT_0 = 16'h0000;
defparam ram16s_inst_17.INIT_1 = 16'h0000;
defparam ram16s_inst_17.INIT_2 = 16'h0000;
defparam ram16s_inst_17.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_18 (
    .DO(ram16s_inst_18_dout[75:72]),
    .DI(di[75:72]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_18.INIT_0 = 16'h0000;
defparam ram16s_inst_18.INIT_1 = 16'h0000;
defparam ram16s_inst_18.INIT_2 = 16'h0000;
defparam ram16s_inst_18.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_19 (
    .DO(ram16s_inst_19_dout[79:76]),
    .DI(di[79:76]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_19.INIT_0 = 16'h0000;
defparam ram16s_inst_19.INIT_1 = 16'h0000;
defparam ram16s_inst_19.INIT_2 = 16'h0000;
defparam ram16s_inst_19.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_20 (
    .DO(ram16s_inst_20_dout[83:80]),
    .DI(di[83:80]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_20.INIT_0 = 16'h0000;
defparam ram16s_inst_20.INIT_1 = 16'h0000;
defparam ram16s_inst_20.INIT_2 = 16'h0000;
defparam ram16s_inst_20.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_21 (
    .DO(ram16s_inst_21_dout[87:84]),
    .DI(di[87:84]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_21.INIT_0 = 16'h0000;
defparam ram16s_inst_21.INIT_1 = 16'h0000;
defparam ram16s_inst_21.INIT_2 = 16'h0000;
defparam ram16s_inst_21.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_22 (
    .DO(ram16s_inst_22_dout[91:88]),
    .DI(di[91:88]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_22.INIT_0 = 16'h0000;
defparam ram16s_inst_22.INIT_1 = 16'h0000;
defparam ram16s_inst_22.INIT_2 = 16'h0000;
defparam ram16s_inst_22.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_23 (
    .DO(ram16s_inst_23_dout[95:92]),
    .DI(di[95:92]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_23.INIT_0 = 16'h0000;
defparam ram16s_inst_23.INIT_1 = 16'h0000;
defparam ram16s_inst_23.INIT_2 = 16'h0000;
defparam ram16s_inst_23.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_24 (
    .DO(ram16s_inst_24_dout[99:96]),
    .DI(di[99:96]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_24.INIT_0 = 16'h0000;
defparam ram16s_inst_24.INIT_1 = 16'h0000;
defparam ram16s_inst_24.INIT_2 = 16'h0000;
defparam ram16s_inst_24.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_25 (
    .DO(ram16s_inst_25_dout[103:100]),
    .DI(di[103:100]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_25.INIT_0 = 16'h0000;
defparam ram16s_inst_25.INIT_1 = 16'h0000;
defparam ram16s_inst_25.INIT_2 = 16'h0000;
defparam ram16s_inst_25.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_26 (
    .DO(ram16s_inst_26_dout[107:104]),
    .DI(di[107:104]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_26.INIT_0 = 16'h0000;
defparam ram16s_inst_26.INIT_1 = 16'h0000;
defparam ram16s_inst_26.INIT_2 = 16'h0000;
defparam ram16s_inst_26.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_27 (
    .DO(ram16s_inst_27_dout[111:108]),
    .DI(di[111:108]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_27.INIT_0 = 16'h0000;
defparam ram16s_inst_27.INIT_1 = 16'h0000;
defparam ram16s_inst_27.INIT_2 = 16'h0000;
defparam ram16s_inst_27.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_28 (
    .DO(ram16s_inst_28_dout[115:112]),
    .DI(di[115:112]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_28.INIT_0 = 16'h0000;
defparam ram16s_inst_28.INIT_1 = 16'h0000;
defparam ram16s_inst_28.INIT_2 = 16'h0000;
defparam ram16s_inst_28.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_29 (
    .DO(ram16s_inst_29_dout[119:116]),
    .DI(di[119:116]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_29.INIT_0 = 16'h0000;
defparam ram16s_inst_29.INIT_1 = 16'h0000;
defparam ram16s_inst_29.INIT_2 = 16'h0000;
defparam ram16s_inst_29.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_30 (
    .DO(ram16s_inst_30_dout[123:120]),
    .DI(di[123:120]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_30.INIT_0 = 16'h0000;
defparam ram16s_inst_30.INIT_1 = 16'h0000;
defparam ram16s_inst_30.INIT_2 = 16'h0000;
defparam ram16s_inst_30.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_31 (
    .DO(ram16s_inst_31_dout[127:124]),
    .DI(di[127:124]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_31.INIT_0 = 16'h0000;
defparam ram16s_inst_31.INIT_1 = 16'h0000;
defparam ram16s_inst_31.INIT_2 = 16'h0000;
defparam ram16s_inst_31.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_32 (
    .DO(ram16s_inst_32_dout[131:128]),
    .DI(di[131:128]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_32.INIT_0 = 16'h0000;
defparam ram16s_inst_32.INIT_1 = 16'h0000;
defparam ram16s_inst_32.INIT_2 = 16'h0000;
defparam ram16s_inst_32.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_33 (
    .DO(ram16s_inst_33_dout[135:132]),
    .DI(di[135:132]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_33.INIT_0 = 16'h0000;
defparam ram16s_inst_33.INIT_1 = 16'h0000;
defparam ram16s_inst_33.INIT_2 = 16'h0000;
defparam ram16s_inst_33.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_34 (
    .DO(ram16s_inst_34_dout[139:136]),
    .DI(di[139:136]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_34.INIT_0 = 16'h0000;
defparam ram16s_inst_34.INIT_1 = 16'h0000;
defparam ram16s_inst_34.INIT_2 = 16'h0000;
defparam ram16s_inst_34.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_35 (
    .DO(ram16s_inst_35_dout[143:140]),
    .DI(di[143:140]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_35.INIT_0 = 16'h0000;
defparam ram16s_inst_35.INIT_1 = 16'h0000;
defparam ram16s_inst_35.INIT_2 = 16'h0000;
defparam ram16s_inst_35.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_36 (
    .DO(ram16s_inst_36_dout[147:144]),
    .DI(di[147:144]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_36.INIT_0 = 16'h0000;
defparam ram16s_inst_36.INIT_1 = 16'h0000;
defparam ram16s_inst_36.INIT_2 = 16'h0000;
defparam ram16s_inst_36.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_37 (
    .DO(ram16s_inst_37_dout[151:148]),
    .DI(di[151:148]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_37.INIT_0 = 16'h0000;
defparam ram16s_inst_37.INIT_1 = 16'h0000;
defparam ram16s_inst_37.INIT_2 = 16'h0000;
defparam ram16s_inst_37.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_38 (
    .DO(ram16s_inst_38_dout[155:152]),
    .DI(di[155:152]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_38.INIT_0 = 16'h0000;
defparam ram16s_inst_38.INIT_1 = 16'h0000;
defparam ram16s_inst_38.INIT_2 = 16'h0000;
defparam ram16s_inst_38.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_39 (
    .DO(ram16s_inst_39_dout[159:156]),
    .DI(di[159:156]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_39.INIT_0 = 16'h0000;
defparam ram16s_inst_39.INIT_1 = 16'h0000;
defparam ram16s_inst_39.INIT_2 = 16'h0000;
defparam ram16s_inst_39.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_40 (
    .DO(ram16s_inst_40_dout[163:160]),
    .DI(di[163:160]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_40.INIT_0 = 16'h0000;
defparam ram16s_inst_40.INIT_1 = 16'h0000;
defparam ram16s_inst_40.INIT_2 = 16'h0000;
defparam ram16s_inst_40.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_41 (
    .DO(ram16s_inst_41_dout[167:164]),
    .DI(di[167:164]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_41.INIT_0 = 16'h0000;
defparam ram16s_inst_41.INIT_1 = 16'h0000;
defparam ram16s_inst_41.INIT_2 = 16'h0000;
defparam ram16s_inst_41.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_42 (
    .DO(ram16s_inst_42_dout[171:168]),
    .DI(di[171:168]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_42.INIT_0 = 16'h0000;
defparam ram16s_inst_42.INIT_1 = 16'h0000;
defparam ram16s_inst_42.INIT_2 = 16'h0000;
defparam ram16s_inst_42.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_43 (
    .DO(ram16s_inst_43_dout[175:172]),
    .DI(di[175:172]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_43.INIT_0 = 16'h0000;
defparam ram16s_inst_43.INIT_1 = 16'h0000;
defparam ram16s_inst_43.INIT_2 = 16'h0000;
defparam ram16s_inst_43.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_44 (
    .DO(ram16s_inst_44_dout[179:176]),
    .DI(di[179:176]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_44.INIT_0 = 16'h0000;
defparam ram16s_inst_44.INIT_1 = 16'h0000;
defparam ram16s_inst_44.INIT_2 = 16'h0000;
defparam ram16s_inst_44.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_45 (
    .DO(ram16s_inst_45_dout[183:180]),
    .DI(di[183:180]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_45.INIT_0 = 16'h0000;
defparam ram16s_inst_45.INIT_1 = 16'h0000;
defparam ram16s_inst_45.INIT_2 = 16'h0000;
defparam ram16s_inst_45.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_46 (
    .DO(ram16s_inst_46_dout[187:184]),
    .DI(di[187:184]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_46.INIT_0 = 16'h0000;
defparam ram16s_inst_46.INIT_1 = 16'h0000;
defparam ram16s_inst_46.INIT_2 = 16'h0000;
defparam ram16s_inst_46.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_47 (
    .DO(ram16s_inst_47_dout[191:188]),
    .DI(di[191:188]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_47.INIT_0 = 16'h0000;
defparam ram16s_inst_47.INIT_1 = 16'h0000;
defparam ram16s_inst_47.INIT_2 = 16'h0000;
defparam ram16s_inst_47.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_48 (
    .DO(ram16s_inst_48_dout[195:192]),
    .DI(di[195:192]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_48.INIT_0 = 16'h0000;
defparam ram16s_inst_48.INIT_1 = 16'h0000;
defparam ram16s_inst_48.INIT_2 = 16'h0000;
defparam ram16s_inst_48.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_49 (
    .DO(ram16s_inst_49_dout[199:196]),
    .DI(di[199:196]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_49.INIT_0 = 16'h0000;
defparam ram16s_inst_49.INIT_1 = 16'h0000;
defparam ram16s_inst_49.INIT_2 = 16'h0000;
defparam ram16s_inst_49.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_50 (
    .DO(ram16s_inst_50_dout[203:200]),
    .DI(di[203:200]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_50.INIT_0 = 16'h0000;
defparam ram16s_inst_50.INIT_1 = 16'h0000;
defparam ram16s_inst_50.INIT_2 = 16'h0000;
defparam ram16s_inst_50.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_51 (
    .DO(ram16s_inst_51_dout[207:204]),
    .DI(di[207:204]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_51.INIT_0 = 16'h0000;
defparam ram16s_inst_51.INIT_1 = 16'h0000;
defparam ram16s_inst_51.INIT_2 = 16'h0000;
defparam ram16s_inst_51.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_52 (
    .DO(ram16s_inst_52_dout[211:208]),
    .DI(di[211:208]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_52.INIT_0 = 16'h0000;
defparam ram16s_inst_52.INIT_1 = 16'h0000;
defparam ram16s_inst_52.INIT_2 = 16'h0000;
defparam ram16s_inst_52.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_53 (
    .DO(ram16s_inst_53_dout[215:212]),
    .DI(di[215:212]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_53.INIT_0 = 16'h0000;
defparam ram16s_inst_53.INIT_1 = 16'h0000;
defparam ram16s_inst_53.INIT_2 = 16'h0000;
defparam ram16s_inst_53.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_54 (
    .DO(ram16s_inst_54_dout[219:216]),
    .DI(di[219:216]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_54.INIT_0 = 16'h0000;
defparam ram16s_inst_54.INIT_1 = 16'h0000;
defparam ram16s_inst_54.INIT_2 = 16'h0000;
defparam ram16s_inst_54.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_55 (
    .DO(ram16s_inst_55_dout[223:220]),
    .DI(di[223:220]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_55.INIT_0 = 16'h0000;
defparam ram16s_inst_55.INIT_1 = 16'h0000;
defparam ram16s_inst_55.INIT_2 = 16'h0000;
defparam ram16s_inst_55.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_56 (
    .DO(ram16s_inst_56_dout[227:224]),
    .DI(di[227:224]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_56.INIT_0 = 16'h0000;
defparam ram16s_inst_56.INIT_1 = 16'h0000;
defparam ram16s_inst_56.INIT_2 = 16'h0000;
defparam ram16s_inst_56.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_57 (
    .DO(ram16s_inst_57_dout[231:228]),
    .DI(di[231:228]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_57.INIT_0 = 16'h0000;
defparam ram16s_inst_57.INIT_1 = 16'h0000;
defparam ram16s_inst_57.INIT_2 = 16'h0000;
defparam ram16s_inst_57.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_58 (
    .DO(ram16s_inst_58_dout[235:232]),
    .DI(di[235:232]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_58.INIT_0 = 16'h0000;
defparam ram16s_inst_58.INIT_1 = 16'h0000;
defparam ram16s_inst_58.INIT_2 = 16'h0000;
defparam ram16s_inst_58.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_59 (
    .DO(ram16s_inst_59_dout[239:236]),
    .DI(di[239:236]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_59.INIT_0 = 16'h0000;
defparam ram16s_inst_59.INIT_1 = 16'h0000;
defparam ram16s_inst_59.INIT_2 = 16'h0000;
defparam ram16s_inst_59.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_60 (
    .DO(ram16s_inst_60_dout[243:240]),
    .DI(di[243:240]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_60.INIT_0 = 16'h0000;
defparam ram16s_inst_60.INIT_1 = 16'h0000;
defparam ram16s_inst_60.INIT_2 = 16'h0000;
defparam ram16s_inst_60.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_61 (
    .DO(ram16s_inst_61_dout[247:244]),
    .DI(di[247:244]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_61.INIT_0 = 16'h0000;
defparam ram16s_inst_61.INIT_1 = 16'h0000;
defparam ram16s_inst_61.INIT_2 = 16'h0000;
defparam ram16s_inst_61.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_62 (
    .DO(ram16s_inst_62_dout[251:248]),
    .DI(di[251:248]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_62.INIT_0 = 16'h0000;
defparam ram16s_inst_62.INIT_1 = 16'h0000;
defparam ram16s_inst_62.INIT_2 = 16'h0000;
defparam ram16s_inst_62.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_63 (
    .DO(ram16s_inst_63_dout[255:252]),
    .DI(di[255:252]),
    .AD(ad[3:0]),
    .WRE(lut_f_0),
    .CLK(clk)
);

defparam ram16s_inst_63.INIT_0 = 16'h0000;
defparam ram16s_inst_63.INIT_1 = 16'h0000;
defparam ram16s_inst_63.INIT_2 = 16'h0000;
defparam ram16s_inst_63.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_64 (
    .DO(ram16s_inst_64_dout[3:0]),
    .DI(di[3:0]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_64.INIT_0 = 16'h0000;
defparam ram16s_inst_64.INIT_1 = 16'h0000;
defparam ram16s_inst_64.INIT_2 = 16'h0000;
defparam ram16s_inst_64.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_65 (
    .DO(ram16s_inst_65_dout[7:4]),
    .DI(di[7:4]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_65.INIT_0 = 16'h0000;
defparam ram16s_inst_65.INIT_1 = 16'h0000;
defparam ram16s_inst_65.INIT_2 = 16'h0000;
defparam ram16s_inst_65.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_66 (
    .DO(ram16s_inst_66_dout[11:8]),
    .DI(di[11:8]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_66.INIT_0 = 16'h0000;
defparam ram16s_inst_66.INIT_1 = 16'h0000;
defparam ram16s_inst_66.INIT_2 = 16'h0000;
defparam ram16s_inst_66.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_67 (
    .DO(ram16s_inst_67_dout[15:12]),
    .DI(di[15:12]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_67.INIT_0 = 16'h0000;
defparam ram16s_inst_67.INIT_1 = 16'h0000;
defparam ram16s_inst_67.INIT_2 = 16'h0000;
defparam ram16s_inst_67.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_68 (
    .DO(ram16s_inst_68_dout[19:16]),
    .DI(di[19:16]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_68.INIT_0 = 16'h0000;
defparam ram16s_inst_68.INIT_1 = 16'h0000;
defparam ram16s_inst_68.INIT_2 = 16'h0000;
defparam ram16s_inst_68.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_69 (
    .DO(ram16s_inst_69_dout[23:20]),
    .DI(di[23:20]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_69.INIT_0 = 16'h0000;
defparam ram16s_inst_69.INIT_1 = 16'h0000;
defparam ram16s_inst_69.INIT_2 = 16'h0000;
defparam ram16s_inst_69.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_70 (
    .DO(ram16s_inst_70_dout[27:24]),
    .DI(di[27:24]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_70.INIT_0 = 16'h0000;
defparam ram16s_inst_70.INIT_1 = 16'h0000;
defparam ram16s_inst_70.INIT_2 = 16'h0000;
defparam ram16s_inst_70.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_71 (
    .DO(ram16s_inst_71_dout[31:28]),
    .DI(di[31:28]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_71.INIT_0 = 16'h0000;
defparam ram16s_inst_71.INIT_1 = 16'h0000;
defparam ram16s_inst_71.INIT_2 = 16'h0000;
defparam ram16s_inst_71.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_72 (
    .DO(ram16s_inst_72_dout[35:32]),
    .DI(di[35:32]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_72.INIT_0 = 16'h0000;
defparam ram16s_inst_72.INIT_1 = 16'h0000;
defparam ram16s_inst_72.INIT_2 = 16'h0000;
defparam ram16s_inst_72.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_73 (
    .DO(ram16s_inst_73_dout[39:36]),
    .DI(di[39:36]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_73.INIT_0 = 16'h0000;
defparam ram16s_inst_73.INIT_1 = 16'h0000;
defparam ram16s_inst_73.INIT_2 = 16'h0000;
defparam ram16s_inst_73.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_74 (
    .DO(ram16s_inst_74_dout[43:40]),
    .DI(di[43:40]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_74.INIT_0 = 16'h0000;
defparam ram16s_inst_74.INIT_1 = 16'h0000;
defparam ram16s_inst_74.INIT_2 = 16'h0000;
defparam ram16s_inst_74.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_75 (
    .DO(ram16s_inst_75_dout[47:44]),
    .DI(di[47:44]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_75.INIT_0 = 16'h0000;
defparam ram16s_inst_75.INIT_1 = 16'h0000;
defparam ram16s_inst_75.INIT_2 = 16'h0000;
defparam ram16s_inst_75.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_76 (
    .DO(ram16s_inst_76_dout[51:48]),
    .DI(di[51:48]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_76.INIT_0 = 16'h0000;
defparam ram16s_inst_76.INIT_1 = 16'h0000;
defparam ram16s_inst_76.INIT_2 = 16'h0000;
defparam ram16s_inst_76.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_77 (
    .DO(ram16s_inst_77_dout[55:52]),
    .DI(di[55:52]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_77.INIT_0 = 16'h0000;
defparam ram16s_inst_77.INIT_1 = 16'h0000;
defparam ram16s_inst_77.INIT_2 = 16'h0000;
defparam ram16s_inst_77.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_78 (
    .DO(ram16s_inst_78_dout[59:56]),
    .DI(di[59:56]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_78.INIT_0 = 16'h0000;
defparam ram16s_inst_78.INIT_1 = 16'h0000;
defparam ram16s_inst_78.INIT_2 = 16'h0000;
defparam ram16s_inst_78.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_79 (
    .DO(ram16s_inst_79_dout[63:60]),
    .DI(di[63:60]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_79.INIT_0 = 16'h0000;
defparam ram16s_inst_79.INIT_1 = 16'h0000;
defparam ram16s_inst_79.INIT_2 = 16'h0000;
defparam ram16s_inst_79.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_80 (
    .DO(ram16s_inst_80_dout[67:64]),
    .DI(di[67:64]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_80.INIT_0 = 16'h0000;
defparam ram16s_inst_80.INIT_1 = 16'h0000;
defparam ram16s_inst_80.INIT_2 = 16'h0000;
defparam ram16s_inst_80.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_81 (
    .DO(ram16s_inst_81_dout[71:68]),
    .DI(di[71:68]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_81.INIT_0 = 16'h0000;
defparam ram16s_inst_81.INIT_1 = 16'h0000;
defparam ram16s_inst_81.INIT_2 = 16'h0000;
defparam ram16s_inst_81.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_82 (
    .DO(ram16s_inst_82_dout[75:72]),
    .DI(di[75:72]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_82.INIT_0 = 16'h0000;
defparam ram16s_inst_82.INIT_1 = 16'h0000;
defparam ram16s_inst_82.INIT_2 = 16'h0000;
defparam ram16s_inst_82.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_83 (
    .DO(ram16s_inst_83_dout[79:76]),
    .DI(di[79:76]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_83.INIT_0 = 16'h0000;
defparam ram16s_inst_83.INIT_1 = 16'h0000;
defparam ram16s_inst_83.INIT_2 = 16'h0000;
defparam ram16s_inst_83.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_84 (
    .DO(ram16s_inst_84_dout[83:80]),
    .DI(di[83:80]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_84.INIT_0 = 16'h0000;
defparam ram16s_inst_84.INIT_1 = 16'h0000;
defparam ram16s_inst_84.INIT_2 = 16'h0000;
defparam ram16s_inst_84.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_85 (
    .DO(ram16s_inst_85_dout[87:84]),
    .DI(di[87:84]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_85.INIT_0 = 16'h0000;
defparam ram16s_inst_85.INIT_1 = 16'h0000;
defparam ram16s_inst_85.INIT_2 = 16'h0000;
defparam ram16s_inst_85.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_86 (
    .DO(ram16s_inst_86_dout[91:88]),
    .DI(di[91:88]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_86.INIT_0 = 16'h0000;
defparam ram16s_inst_86.INIT_1 = 16'h0000;
defparam ram16s_inst_86.INIT_2 = 16'h0000;
defparam ram16s_inst_86.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_87 (
    .DO(ram16s_inst_87_dout[95:92]),
    .DI(di[95:92]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_87.INIT_0 = 16'h0000;
defparam ram16s_inst_87.INIT_1 = 16'h0000;
defparam ram16s_inst_87.INIT_2 = 16'h0000;
defparam ram16s_inst_87.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_88 (
    .DO(ram16s_inst_88_dout[99:96]),
    .DI(di[99:96]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_88.INIT_0 = 16'h0000;
defparam ram16s_inst_88.INIT_1 = 16'h0000;
defparam ram16s_inst_88.INIT_2 = 16'h0000;
defparam ram16s_inst_88.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_89 (
    .DO(ram16s_inst_89_dout[103:100]),
    .DI(di[103:100]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_89.INIT_0 = 16'h0000;
defparam ram16s_inst_89.INIT_1 = 16'h0000;
defparam ram16s_inst_89.INIT_2 = 16'h0000;
defparam ram16s_inst_89.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_90 (
    .DO(ram16s_inst_90_dout[107:104]),
    .DI(di[107:104]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_90.INIT_0 = 16'h0000;
defparam ram16s_inst_90.INIT_1 = 16'h0000;
defparam ram16s_inst_90.INIT_2 = 16'h0000;
defparam ram16s_inst_90.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_91 (
    .DO(ram16s_inst_91_dout[111:108]),
    .DI(di[111:108]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_91.INIT_0 = 16'h0000;
defparam ram16s_inst_91.INIT_1 = 16'h0000;
defparam ram16s_inst_91.INIT_2 = 16'h0000;
defparam ram16s_inst_91.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_92 (
    .DO(ram16s_inst_92_dout[115:112]),
    .DI(di[115:112]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_92.INIT_0 = 16'h0000;
defparam ram16s_inst_92.INIT_1 = 16'h0000;
defparam ram16s_inst_92.INIT_2 = 16'h0000;
defparam ram16s_inst_92.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_93 (
    .DO(ram16s_inst_93_dout[119:116]),
    .DI(di[119:116]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_93.INIT_0 = 16'h0000;
defparam ram16s_inst_93.INIT_1 = 16'h0000;
defparam ram16s_inst_93.INIT_2 = 16'h0000;
defparam ram16s_inst_93.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_94 (
    .DO(ram16s_inst_94_dout[123:120]),
    .DI(di[123:120]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_94.INIT_0 = 16'h0000;
defparam ram16s_inst_94.INIT_1 = 16'h0000;
defparam ram16s_inst_94.INIT_2 = 16'h0000;
defparam ram16s_inst_94.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_95 (
    .DO(ram16s_inst_95_dout[127:124]),
    .DI(di[127:124]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_95.INIT_0 = 16'h0000;
defparam ram16s_inst_95.INIT_1 = 16'h0000;
defparam ram16s_inst_95.INIT_2 = 16'h0000;
defparam ram16s_inst_95.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_96 (
    .DO(ram16s_inst_96_dout[131:128]),
    .DI(di[131:128]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_96.INIT_0 = 16'h0000;
defparam ram16s_inst_96.INIT_1 = 16'h0000;
defparam ram16s_inst_96.INIT_2 = 16'h0000;
defparam ram16s_inst_96.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_97 (
    .DO(ram16s_inst_97_dout[135:132]),
    .DI(di[135:132]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_97.INIT_0 = 16'h0000;
defparam ram16s_inst_97.INIT_1 = 16'h0000;
defparam ram16s_inst_97.INIT_2 = 16'h0000;
defparam ram16s_inst_97.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_98 (
    .DO(ram16s_inst_98_dout[139:136]),
    .DI(di[139:136]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_98.INIT_0 = 16'h0000;
defparam ram16s_inst_98.INIT_1 = 16'h0000;
defparam ram16s_inst_98.INIT_2 = 16'h0000;
defparam ram16s_inst_98.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_99 (
    .DO(ram16s_inst_99_dout[143:140]),
    .DI(di[143:140]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_99.INIT_0 = 16'h0000;
defparam ram16s_inst_99.INIT_1 = 16'h0000;
defparam ram16s_inst_99.INIT_2 = 16'h0000;
defparam ram16s_inst_99.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_100 (
    .DO(ram16s_inst_100_dout[147:144]),
    .DI(di[147:144]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_100.INIT_0 = 16'h0000;
defparam ram16s_inst_100.INIT_1 = 16'h0000;
defparam ram16s_inst_100.INIT_2 = 16'h0000;
defparam ram16s_inst_100.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_101 (
    .DO(ram16s_inst_101_dout[151:148]),
    .DI(di[151:148]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_101.INIT_0 = 16'h0000;
defparam ram16s_inst_101.INIT_1 = 16'h0000;
defparam ram16s_inst_101.INIT_2 = 16'h0000;
defparam ram16s_inst_101.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_102 (
    .DO(ram16s_inst_102_dout[155:152]),
    .DI(di[155:152]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_102.INIT_0 = 16'h0000;
defparam ram16s_inst_102.INIT_1 = 16'h0000;
defparam ram16s_inst_102.INIT_2 = 16'h0000;
defparam ram16s_inst_102.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_103 (
    .DO(ram16s_inst_103_dout[159:156]),
    .DI(di[159:156]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_103.INIT_0 = 16'h0000;
defparam ram16s_inst_103.INIT_1 = 16'h0000;
defparam ram16s_inst_103.INIT_2 = 16'h0000;
defparam ram16s_inst_103.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_104 (
    .DO(ram16s_inst_104_dout[163:160]),
    .DI(di[163:160]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_104.INIT_0 = 16'h0000;
defparam ram16s_inst_104.INIT_1 = 16'h0000;
defparam ram16s_inst_104.INIT_2 = 16'h0000;
defparam ram16s_inst_104.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_105 (
    .DO(ram16s_inst_105_dout[167:164]),
    .DI(di[167:164]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_105.INIT_0 = 16'h0000;
defparam ram16s_inst_105.INIT_1 = 16'h0000;
defparam ram16s_inst_105.INIT_2 = 16'h0000;
defparam ram16s_inst_105.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_106 (
    .DO(ram16s_inst_106_dout[171:168]),
    .DI(di[171:168]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_106.INIT_0 = 16'h0000;
defparam ram16s_inst_106.INIT_1 = 16'h0000;
defparam ram16s_inst_106.INIT_2 = 16'h0000;
defparam ram16s_inst_106.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_107 (
    .DO(ram16s_inst_107_dout[175:172]),
    .DI(di[175:172]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_107.INIT_0 = 16'h0000;
defparam ram16s_inst_107.INIT_1 = 16'h0000;
defparam ram16s_inst_107.INIT_2 = 16'h0000;
defparam ram16s_inst_107.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_108 (
    .DO(ram16s_inst_108_dout[179:176]),
    .DI(di[179:176]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_108.INIT_0 = 16'h0000;
defparam ram16s_inst_108.INIT_1 = 16'h0000;
defparam ram16s_inst_108.INIT_2 = 16'h0000;
defparam ram16s_inst_108.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_109 (
    .DO(ram16s_inst_109_dout[183:180]),
    .DI(di[183:180]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_109.INIT_0 = 16'h0000;
defparam ram16s_inst_109.INIT_1 = 16'h0000;
defparam ram16s_inst_109.INIT_2 = 16'h0000;
defparam ram16s_inst_109.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_110 (
    .DO(ram16s_inst_110_dout[187:184]),
    .DI(di[187:184]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_110.INIT_0 = 16'h0000;
defparam ram16s_inst_110.INIT_1 = 16'h0000;
defparam ram16s_inst_110.INIT_2 = 16'h0000;
defparam ram16s_inst_110.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_111 (
    .DO(ram16s_inst_111_dout[191:188]),
    .DI(di[191:188]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_111.INIT_0 = 16'h0000;
defparam ram16s_inst_111.INIT_1 = 16'h0000;
defparam ram16s_inst_111.INIT_2 = 16'h0000;
defparam ram16s_inst_111.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_112 (
    .DO(ram16s_inst_112_dout[195:192]),
    .DI(di[195:192]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_112.INIT_0 = 16'h0000;
defparam ram16s_inst_112.INIT_1 = 16'h0000;
defparam ram16s_inst_112.INIT_2 = 16'h0000;
defparam ram16s_inst_112.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_113 (
    .DO(ram16s_inst_113_dout[199:196]),
    .DI(di[199:196]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_113.INIT_0 = 16'h0000;
defparam ram16s_inst_113.INIT_1 = 16'h0000;
defparam ram16s_inst_113.INIT_2 = 16'h0000;
defparam ram16s_inst_113.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_114 (
    .DO(ram16s_inst_114_dout[203:200]),
    .DI(di[203:200]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_114.INIT_0 = 16'h0000;
defparam ram16s_inst_114.INIT_1 = 16'h0000;
defparam ram16s_inst_114.INIT_2 = 16'h0000;
defparam ram16s_inst_114.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_115 (
    .DO(ram16s_inst_115_dout[207:204]),
    .DI(di[207:204]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_115.INIT_0 = 16'h0000;
defparam ram16s_inst_115.INIT_1 = 16'h0000;
defparam ram16s_inst_115.INIT_2 = 16'h0000;
defparam ram16s_inst_115.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_116 (
    .DO(ram16s_inst_116_dout[211:208]),
    .DI(di[211:208]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_116.INIT_0 = 16'h0000;
defparam ram16s_inst_116.INIT_1 = 16'h0000;
defparam ram16s_inst_116.INIT_2 = 16'h0000;
defparam ram16s_inst_116.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_117 (
    .DO(ram16s_inst_117_dout[215:212]),
    .DI(di[215:212]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_117.INIT_0 = 16'h0000;
defparam ram16s_inst_117.INIT_1 = 16'h0000;
defparam ram16s_inst_117.INIT_2 = 16'h0000;
defparam ram16s_inst_117.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_118 (
    .DO(ram16s_inst_118_dout[219:216]),
    .DI(di[219:216]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_118.INIT_0 = 16'h0000;
defparam ram16s_inst_118.INIT_1 = 16'h0000;
defparam ram16s_inst_118.INIT_2 = 16'h0000;
defparam ram16s_inst_118.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_119 (
    .DO(ram16s_inst_119_dout[223:220]),
    .DI(di[223:220]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_119.INIT_0 = 16'h0000;
defparam ram16s_inst_119.INIT_1 = 16'h0000;
defparam ram16s_inst_119.INIT_2 = 16'h0000;
defparam ram16s_inst_119.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_120 (
    .DO(ram16s_inst_120_dout[227:224]),
    .DI(di[227:224]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_120.INIT_0 = 16'h0000;
defparam ram16s_inst_120.INIT_1 = 16'h0000;
defparam ram16s_inst_120.INIT_2 = 16'h0000;
defparam ram16s_inst_120.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_121 (
    .DO(ram16s_inst_121_dout[231:228]),
    .DI(di[231:228]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_121.INIT_0 = 16'h0000;
defparam ram16s_inst_121.INIT_1 = 16'h0000;
defparam ram16s_inst_121.INIT_2 = 16'h0000;
defparam ram16s_inst_121.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_122 (
    .DO(ram16s_inst_122_dout[235:232]),
    .DI(di[235:232]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_122.INIT_0 = 16'h0000;
defparam ram16s_inst_122.INIT_1 = 16'h0000;
defparam ram16s_inst_122.INIT_2 = 16'h0000;
defparam ram16s_inst_122.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_123 (
    .DO(ram16s_inst_123_dout[239:236]),
    .DI(di[239:236]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_123.INIT_0 = 16'h0000;
defparam ram16s_inst_123.INIT_1 = 16'h0000;
defparam ram16s_inst_123.INIT_2 = 16'h0000;
defparam ram16s_inst_123.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_124 (
    .DO(ram16s_inst_124_dout[243:240]),
    .DI(di[243:240]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_124.INIT_0 = 16'h0000;
defparam ram16s_inst_124.INIT_1 = 16'h0000;
defparam ram16s_inst_124.INIT_2 = 16'h0000;
defparam ram16s_inst_124.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_125 (
    .DO(ram16s_inst_125_dout[247:244]),
    .DI(di[247:244]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_125.INIT_0 = 16'h0000;
defparam ram16s_inst_125.INIT_1 = 16'h0000;
defparam ram16s_inst_125.INIT_2 = 16'h0000;
defparam ram16s_inst_125.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_126 (
    .DO(ram16s_inst_126_dout[251:248]),
    .DI(di[251:248]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_126.INIT_0 = 16'h0000;
defparam ram16s_inst_126.INIT_1 = 16'h0000;
defparam ram16s_inst_126.INIT_2 = 16'h0000;
defparam ram16s_inst_126.INIT_3 = 16'h0000;

RAM16S4 ram16s_inst_127 (
    .DO(ram16s_inst_127_dout[255:252]),
    .DI(di[255:252]),
    .AD(ad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16s_inst_127.INIT_0 = 16'h0000;
defparam ram16s_inst_127.INIT_1 = 16'h0000;
defparam ram16s_inst_127.INIT_2 = 16'h0000;
defparam ram16s_inst_127.INIT_3 = 16'h0000;

MUX2 mux_inst_0 (
  .O(dout[0]),
  .I0(ram16s_inst_0_dout[0]),
  .I1(ram16s_inst_64_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_1 (
  .O(dout[1]),
  .I0(ram16s_inst_0_dout[1]),
  .I1(ram16s_inst_64_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_2 (
  .O(dout[2]),
  .I0(ram16s_inst_0_dout[2]),
  .I1(ram16s_inst_64_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_3 (
  .O(dout[3]),
  .I0(ram16s_inst_0_dout[3]),
  .I1(ram16s_inst_64_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_4 (
  .O(dout[4]),
  .I0(ram16s_inst_1_dout[4]),
  .I1(ram16s_inst_65_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_5 (
  .O(dout[5]),
  .I0(ram16s_inst_1_dout[5]),
  .I1(ram16s_inst_65_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_6 (
  .O(dout[6]),
  .I0(ram16s_inst_1_dout[6]),
  .I1(ram16s_inst_65_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_7 (
  .O(dout[7]),
  .I0(ram16s_inst_1_dout[7]),
  .I1(ram16s_inst_65_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_8 (
  .O(dout[8]),
  .I0(ram16s_inst_2_dout[8]),
  .I1(ram16s_inst_66_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_9 (
  .O(dout[9]),
  .I0(ram16s_inst_2_dout[9]),
  .I1(ram16s_inst_66_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_10 (
  .O(dout[10]),
  .I0(ram16s_inst_2_dout[10]),
  .I1(ram16s_inst_66_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_11 (
  .O(dout[11]),
  .I0(ram16s_inst_2_dout[11]),
  .I1(ram16s_inst_66_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_12 (
  .O(dout[12]),
  .I0(ram16s_inst_3_dout[12]),
  .I1(ram16s_inst_67_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_13 (
  .O(dout[13]),
  .I0(ram16s_inst_3_dout[13]),
  .I1(ram16s_inst_67_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_14 (
  .O(dout[14]),
  .I0(ram16s_inst_3_dout[14]),
  .I1(ram16s_inst_67_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_15 (
  .O(dout[15]),
  .I0(ram16s_inst_3_dout[15]),
  .I1(ram16s_inst_67_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_16 (
  .O(dout[16]),
  .I0(ram16s_inst_4_dout[16]),
  .I1(ram16s_inst_68_dout[16]),
  .S0(ad[4])
);
MUX2 mux_inst_17 (
  .O(dout[17]),
  .I0(ram16s_inst_4_dout[17]),
  .I1(ram16s_inst_68_dout[17]),
  .S0(ad[4])
);
MUX2 mux_inst_18 (
  .O(dout[18]),
  .I0(ram16s_inst_4_dout[18]),
  .I1(ram16s_inst_68_dout[18]),
  .S0(ad[4])
);
MUX2 mux_inst_19 (
  .O(dout[19]),
  .I0(ram16s_inst_4_dout[19]),
  .I1(ram16s_inst_68_dout[19]),
  .S0(ad[4])
);
MUX2 mux_inst_20 (
  .O(dout[20]),
  .I0(ram16s_inst_5_dout[20]),
  .I1(ram16s_inst_69_dout[20]),
  .S0(ad[4])
);
MUX2 mux_inst_21 (
  .O(dout[21]),
  .I0(ram16s_inst_5_dout[21]),
  .I1(ram16s_inst_69_dout[21]),
  .S0(ad[4])
);
MUX2 mux_inst_22 (
  .O(dout[22]),
  .I0(ram16s_inst_5_dout[22]),
  .I1(ram16s_inst_69_dout[22]),
  .S0(ad[4])
);
MUX2 mux_inst_23 (
  .O(dout[23]),
  .I0(ram16s_inst_5_dout[23]),
  .I1(ram16s_inst_69_dout[23]),
  .S0(ad[4])
);
MUX2 mux_inst_24 (
  .O(dout[24]),
  .I0(ram16s_inst_6_dout[24]),
  .I1(ram16s_inst_70_dout[24]),
  .S0(ad[4])
);
MUX2 mux_inst_25 (
  .O(dout[25]),
  .I0(ram16s_inst_6_dout[25]),
  .I1(ram16s_inst_70_dout[25]),
  .S0(ad[4])
);
MUX2 mux_inst_26 (
  .O(dout[26]),
  .I0(ram16s_inst_6_dout[26]),
  .I1(ram16s_inst_70_dout[26]),
  .S0(ad[4])
);
MUX2 mux_inst_27 (
  .O(dout[27]),
  .I0(ram16s_inst_6_dout[27]),
  .I1(ram16s_inst_70_dout[27]),
  .S0(ad[4])
);
MUX2 mux_inst_28 (
  .O(dout[28]),
  .I0(ram16s_inst_7_dout[28]),
  .I1(ram16s_inst_71_dout[28]),
  .S0(ad[4])
);
MUX2 mux_inst_29 (
  .O(dout[29]),
  .I0(ram16s_inst_7_dout[29]),
  .I1(ram16s_inst_71_dout[29]),
  .S0(ad[4])
);
MUX2 mux_inst_30 (
  .O(dout[30]),
  .I0(ram16s_inst_7_dout[30]),
  .I1(ram16s_inst_71_dout[30]),
  .S0(ad[4])
);
MUX2 mux_inst_31 (
  .O(dout[31]),
  .I0(ram16s_inst_7_dout[31]),
  .I1(ram16s_inst_71_dout[31]),
  .S0(ad[4])
);
MUX2 mux_inst_32 (
  .O(dout[32]),
  .I0(ram16s_inst_8_dout[32]),
  .I1(ram16s_inst_72_dout[32]),
  .S0(ad[4])
);
MUX2 mux_inst_33 (
  .O(dout[33]),
  .I0(ram16s_inst_8_dout[33]),
  .I1(ram16s_inst_72_dout[33]),
  .S0(ad[4])
);
MUX2 mux_inst_34 (
  .O(dout[34]),
  .I0(ram16s_inst_8_dout[34]),
  .I1(ram16s_inst_72_dout[34]),
  .S0(ad[4])
);
MUX2 mux_inst_35 (
  .O(dout[35]),
  .I0(ram16s_inst_8_dout[35]),
  .I1(ram16s_inst_72_dout[35]),
  .S0(ad[4])
);
MUX2 mux_inst_36 (
  .O(dout[36]),
  .I0(ram16s_inst_9_dout[36]),
  .I1(ram16s_inst_73_dout[36]),
  .S0(ad[4])
);
MUX2 mux_inst_37 (
  .O(dout[37]),
  .I0(ram16s_inst_9_dout[37]),
  .I1(ram16s_inst_73_dout[37]),
  .S0(ad[4])
);
MUX2 mux_inst_38 (
  .O(dout[38]),
  .I0(ram16s_inst_9_dout[38]),
  .I1(ram16s_inst_73_dout[38]),
  .S0(ad[4])
);
MUX2 mux_inst_39 (
  .O(dout[39]),
  .I0(ram16s_inst_9_dout[39]),
  .I1(ram16s_inst_73_dout[39]),
  .S0(ad[4])
);
MUX2 mux_inst_40 (
  .O(dout[40]),
  .I0(ram16s_inst_10_dout[40]),
  .I1(ram16s_inst_74_dout[40]),
  .S0(ad[4])
);
MUX2 mux_inst_41 (
  .O(dout[41]),
  .I0(ram16s_inst_10_dout[41]),
  .I1(ram16s_inst_74_dout[41]),
  .S0(ad[4])
);
MUX2 mux_inst_42 (
  .O(dout[42]),
  .I0(ram16s_inst_10_dout[42]),
  .I1(ram16s_inst_74_dout[42]),
  .S0(ad[4])
);
MUX2 mux_inst_43 (
  .O(dout[43]),
  .I0(ram16s_inst_10_dout[43]),
  .I1(ram16s_inst_74_dout[43]),
  .S0(ad[4])
);
MUX2 mux_inst_44 (
  .O(dout[44]),
  .I0(ram16s_inst_11_dout[44]),
  .I1(ram16s_inst_75_dout[44]),
  .S0(ad[4])
);
MUX2 mux_inst_45 (
  .O(dout[45]),
  .I0(ram16s_inst_11_dout[45]),
  .I1(ram16s_inst_75_dout[45]),
  .S0(ad[4])
);
MUX2 mux_inst_46 (
  .O(dout[46]),
  .I0(ram16s_inst_11_dout[46]),
  .I1(ram16s_inst_75_dout[46]),
  .S0(ad[4])
);
MUX2 mux_inst_47 (
  .O(dout[47]),
  .I0(ram16s_inst_11_dout[47]),
  .I1(ram16s_inst_75_dout[47]),
  .S0(ad[4])
);
MUX2 mux_inst_48 (
  .O(dout[48]),
  .I0(ram16s_inst_12_dout[48]),
  .I1(ram16s_inst_76_dout[48]),
  .S0(ad[4])
);
MUX2 mux_inst_49 (
  .O(dout[49]),
  .I0(ram16s_inst_12_dout[49]),
  .I1(ram16s_inst_76_dout[49]),
  .S0(ad[4])
);
MUX2 mux_inst_50 (
  .O(dout[50]),
  .I0(ram16s_inst_12_dout[50]),
  .I1(ram16s_inst_76_dout[50]),
  .S0(ad[4])
);
MUX2 mux_inst_51 (
  .O(dout[51]),
  .I0(ram16s_inst_12_dout[51]),
  .I1(ram16s_inst_76_dout[51]),
  .S0(ad[4])
);
MUX2 mux_inst_52 (
  .O(dout[52]),
  .I0(ram16s_inst_13_dout[52]),
  .I1(ram16s_inst_77_dout[52]),
  .S0(ad[4])
);
MUX2 mux_inst_53 (
  .O(dout[53]),
  .I0(ram16s_inst_13_dout[53]),
  .I1(ram16s_inst_77_dout[53]),
  .S0(ad[4])
);
MUX2 mux_inst_54 (
  .O(dout[54]),
  .I0(ram16s_inst_13_dout[54]),
  .I1(ram16s_inst_77_dout[54]),
  .S0(ad[4])
);
MUX2 mux_inst_55 (
  .O(dout[55]),
  .I0(ram16s_inst_13_dout[55]),
  .I1(ram16s_inst_77_dout[55]),
  .S0(ad[4])
);
MUX2 mux_inst_56 (
  .O(dout[56]),
  .I0(ram16s_inst_14_dout[56]),
  .I1(ram16s_inst_78_dout[56]),
  .S0(ad[4])
);
MUX2 mux_inst_57 (
  .O(dout[57]),
  .I0(ram16s_inst_14_dout[57]),
  .I1(ram16s_inst_78_dout[57]),
  .S0(ad[4])
);
MUX2 mux_inst_58 (
  .O(dout[58]),
  .I0(ram16s_inst_14_dout[58]),
  .I1(ram16s_inst_78_dout[58]),
  .S0(ad[4])
);
MUX2 mux_inst_59 (
  .O(dout[59]),
  .I0(ram16s_inst_14_dout[59]),
  .I1(ram16s_inst_78_dout[59]),
  .S0(ad[4])
);
MUX2 mux_inst_60 (
  .O(dout[60]),
  .I0(ram16s_inst_15_dout[60]),
  .I1(ram16s_inst_79_dout[60]),
  .S0(ad[4])
);
MUX2 mux_inst_61 (
  .O(dout[61]),
  .I0(ram16s_inst_15_dout[61]),
  .I1(ram16s_inst_79_dout[61]),
  .S0(ad[4])
);
MUX2 mux_inst_62 (
  .O(dout[62]),
  .I0(ram16s_inst_15_dout[62]),
  .I1(ram16s_inst_79_dout[62]),
  .S0(ad[4])
);
MUX2 mux_inst_63 (
  .O(dout[63]),
  .I0(ram16s_inst_15_dout[63]),
  .I1(ram16s_inst_79_dout[63]),
  .S0(ad[4])
);
MUX2 mux_inst_64 (
  .O(dout[64]),
  .I0(ram16s_inst_16_dout[64]),
  .I1(ram16s_inst_80_dout[64]),
  .S0(ad[4])
);
MUX2 mux_inst_65 (
  .O(dout[65]),
  .I0(ram16s_inst_16_dout[65]),
  .I1(ram16s_inst_80_dout[65]),
  .S0(ad[4])
);
MUX2 mux_inst_66 (
  .O(dout[66]),
  .I0(ram16s_inst_16_dout[66]),
  .I1(ram16s_inst_80_dout[66]),
  .S0(ad[4])
);
MUX2 mux_inst_67 (
  .O(dout[67]),
  .I0(ram16s_inst_16_dout[67]),
  .I1(ram16s_inst_80_dout[67]),
  .S0(ad[4])
);
MUX2 mux_inst_68 (
  .O(dout[68]),
  .I0(ram16s_inst_17_dout[68]),
  .I1(ram16s_inst_81_dout[68]),
  .S0(ad[4])
);
MUX2 mux_inst_69 (
  .O(dout[69]),
  .I0(ram16s_inst_17_dout[69]),
  .I1(ram16s_inst_81_dout[69]),
  .S0(ad[4])
);
MUX2 mux_inst_70 (
  .O(dout[70]),
  .I0(ram16s_inst_17_dout[70]),
  .I1(ram16s_inst_81_dout[70]),
  .S0(ad[4])
);
MUX2 mux_inst_71 (
  .O(dout[71]),
  .I0(ram16s_inst_17_dout[71]),
  .I1(ram16s_inst_81_dout[71]),
  .S0(ad[4])
);
MUX2 mux_inst_72 (
  .O(dout[72]),
  .I0(ram16s_inst_18_dout[72]),
  .I1(ram16s_inst_82_dout[72]),
  .S0(ad[4])
);
MUX2 mux_inst_73 (
  .O(dout[73]),
  .I0(ram16s_inst_18_dout[73]),
  .I1(ram16s_inst_82_dout[73]),
  .S0(ad[4])
);
MUX2 mux_inst_74 (
  .O(dout[74]),
  .I0(ram16s_inst_18_dout[74]),
  .I1(ram16s_inst_82_dout[74]),
  .S0(ad[4])
);
MUX2 mux_inst_75 (
  .O(dout[75]),
  .I0(ram16s_inst_18_dout[75]),
  .I1(ram16s_inst_82_dout[75]),
  .S0(ad[4])
);
MUX2 mux_inst_76 (
  .O(dout[76]),
  .I0(ram16s_inst_19_dout[76]),
  .I1(ram16s_inst_83_dout[76]),
  .S0(ad[4])
);
MUX2 mux_inst_77 (
  .O(dout[77]),
  .I0(ram16s_inst_19_dout[77]),
  .I1(ram16s_inst_83_dout[77]),
  .S0(ad[4])
);
MUX2 mux_inst_78 (
  .O(dout[78]),
  .I0(ram16s_inst_19_dout[78]),
  .I1(ram16s_inst_83_dout[78]),
  .S0(ad[4])
);
MUX2 mux_inst_79 (
  .O(dout[79]),
  .I0(ram16s_inst_19_dout[79]),
  .I1(ram16s_inst_83_dout[79]),
  .S0(ad[4])
);
MUX2 mux_inst_80 (
  .O(dout[80]),
  .I0(ram16s_inst_20_dout[80]),
  .I1(ram16s_inst_84_dout[80]),
  .S0(ad[4])
);
MUX2 mux_inst_81 (
  .O(dout[81]),
  .I0(ram16s_inst_20_dout[81]),
  .I1(ram16s_inst_84_dout[81]),
  .S0(ad[4])
);
MUX2 mux_inst_82 (
  .O(dout[82]),
  .I0(ram16s_inst_20_dout[82]),
  .I1(ram16s_inst_84_dout[82]),
  .S0(ad[4])
);
MUX2 mux_inst_83 (
  .O(dout[83]),
  .I0(ram16s_inst_20_dout[83]),
  .I1(ram16s_inst_84_dout[83]),
  .S0(ad[4])
);
MUX2 mux_inst_84 (
  .O(dout[84]),
  .I0(ram16s_inst_21_dout[84]),
  .I1(ram16s_inst_85_dout[84]),
  .S0(ad[4])
);
MUX2 mux_inst_85 (
  .O(dout[85]),
  .I0(ram16s_inst_21_dout[85]),
  .I1(ram16s_inst_85_dout[85]),
  .S0(ad[4])
);
MUX2 mux_inst_86 (
  .O(dout[86]),
  .I0(ram16s_inst_21_dout[86]),
  .I1(ram16s_inst_85_dout[86]),
  .S0(ad[4])
);
MUX2 mux_inst_87 (
  .O(dout[87]),
  .I0(ram16s_inst_21_dout[87]),
  .I1(ram16s_inst_85_dout[87]),
  .S0(ad[4])
);
MUX2 mux_inst_88 (
  .O(dout[88]),
  .I0(ram16s_inst_22_dout[88]),
  .I1(ram16s_inst_86_dout[88]),
  .S0(ad[4])
);
MUX2 mux_inst_89 (
  .O(dout[89]),
  .I0(ram16s_inst_22_dout[89]),
  .I1(ram16s_inst_86_dout[89]),
  .S0(ad[4])
);
MUX2 mux_inst_90 (
  .O(dout[90]),
  .I0(ram16s_inst_22_dout[90]),
  .I1(ram16s_inst_86_dout[90]),
  .S0(ad[4])
);
MUX2 mux_inst_91 (
  .O(dout[91]),
  .I0(ram16s_inst_22_dout[91]),
  .I1(ram16s_inst_86_dout[91]),
  .S0(ad[4])
);
MUX2 mux_inst_92 (
  .O(dout[92]),
  .I0(ram16s_inst_23_dout[92]),
  .I1(ram16s_inst_87_dout[92]),
  .S0(ad[4])
);
MUX2 mux_inst_93 (
  .O(dout[93]),
  .I0(ram16s_inst_23_dout[93]),
  .I1(ram16s_inst_87_dout[93]),
  .S0(ad[4])
);
MUX2 mux_inst_94 (
  .O(dout[94]),
  .I0(ram16s_inst_23_dout[94]),
  .I1(ram16s_inst_87_dout[94]),
  .S0(ad[4])
);
MUX2 mux_inst_95 (
  .O(dout[95]),
  .I0(ram16s_inst_23_dout[95]),
  .I1(ram16s_inst_87_dout[95]),
  .S0(ad[4])
);
MUX2 mux_inst_96 (
  .O(dout[96]),
  .I0(ram16s_inst_24_dout[96]),
  .I1(ram16s_inst_88_dout[96]),
  .S0(ad[4])
);
MUX2 mux_inst_97 (
  .O(dout[97]),
  .I0(ram16s_inst_24_dout[97]),
  .I1(ram16s_inst_88_dout[97]),
  .S0(ad[4])
);
MUX2 mux_inst_98 (
  .O(dout[98]),
  .I0(ram16s_inst_24_dout[98]),
  .I1(ram16s_inst_88_dout[98]),
  .S0(ad[4])
);
MUX2 mux_inst_99 (
  .O(dout[99]),
  .I0(ram16s_inst_24_dout[99]),
  .I1(ram16s_inst_88_dout[99]),
  .S0(ad[4])
);
MUX2 mux_inst_100 (
  .O(dout[100]),
  .I0(ram16s_inst_25_dout[100]),
  .I1(ram16s_inst_89_dout[100]),
  .S0(ad[4])
);
MUX2 mux_inst_101 (
  .O(dout[101]),
  .I0(ram16s_inst_25_dout[101]),
  .I1(ram16s_inst_89_dout[101]),
  .S0(ad[4])
);
MUX2 mux_inst_102 (
  .O(dout[102]),
  .I0(ram16s_inst_25_dout[102]),
  .I1(ram16s_inst_89_dout[102]),
  .S0(ad[4])
);
MUX2 mux_inst_103 (
  .O(dout[103]),
  .I0(ram16s_inst_25_dout[103]),
  .I1(ram16s_inst_89_dout[103]),
  .S0(ad[4])
);
MUX2 mux_inst_104 (
  .O(dout[104]),
  .I0(ram16s_inst_26_dout[104]),
  .I1(ram16s_inst_90_dout[104]),
  .S0(ad[4])
);
MUX2 mux_inst_105 (
  .O(dout[105]),
  .I0(ram16s_inst_26_dout[105]),
  .I1(ram16s_inst_90_dout[105]),
  .S0(ad[4])
);
MUX2 mux_inst_106 (
  .O(dout[106]),
  .I0(ram16s_inst_26_dout[106]),
  .I1(ram16s_inst_90_dout[106]),
  .S0(ad[4])
);
MUX2 mux_inst_107 (
  .O(dout[107]),
  .I0(ram16s_inst_26_dout[107]),
  .I1(ram16s_inst_90_dout[107]),
  .S0(ad[4])
);
MUX2 mux_inst_108 (
  .O(dout[108]),
  .I0(ram16s_inst_27_dout[108]),
  .I1(ram16s_inst_91_dout[108]),
  .S0(ad[4])
);
MUX2 mux_inst_109 (
  .O(dout[109]),
  .I0(ram16s_inst_27_dout[109]),
  .I1(ram16s_inst_91_dout[109]),
  .S0(ad[4])
);
MUX2 mux_inst_110 (
  .O(dout[110]),
  .I0(ram16s_inst_27_dout[110]),
  .I1(ram16s_inst_91_dout[110]),
  .S0(ad[4])
);
MUX2 mux_inst_111 (
  .O(dout[111]),
  .I0(ram16s_inst_27_dout[111]),
  .I1(ram16s_inst_91_dout[111]),
  .S0(ad[4])
);
MUX2 mux_inst_112 (
  .O(dout[112]),
  .I0(ram16s_inst_28_dout[112]),
  .I1(ram16s_inst_92_dout[112]),
  .S0(ad[4])
);
MUX2 mux_inst_113 (
  .O(dout[113]),
  .I0(ram16s_inst_28_dout[113]),
  .I1(ram16s_inst_92_dout[113]),
  .S0(ad[4])
);
MUX2 mux_inst_114 (
  .O(dout[114]),
  .I0(ram16s_inst_28_dout[114]),
  .I1(ram16s_inst_92_dout[114]),
  .S0(ad[4])
);
MUX2 mux_inst_115 (
  .O(dout[115]),
  .I0(ram16s_inst_28_dout[115]),
  .I1(ram16s_inst_92_dout[115]),
  .S0(ad[4])
);
MUX2 mux_inst_116 (
  .O(dout[116]),
  .I0(ram16s_inst_29_dout[116]),
  .I1(ram16s_inst_93_dout[116]),
  .S0(ad[4])
);
MUX2 mux_inst_117 (
  .O(dout[117]),
  .I0(ram16s_inst_29_dout[117]),
  .I1(ram16s_inst_93_dout[117]),
  .S0(ad[4])
);
MUX2 mux_inst_118 (
  .O(dout[118]),
  .I0(ram16s_inst_29_dout[118]),
  .I1(ram16s_inst_93_dout[118]),
  .S0(ad[4])
);
MUX2 mux_inst_119 (
  .O(dout[119]),
  .I0(ram16s_inst_29_dout[119]),
  .I1(ram16s_inst_93_dout[119]),
  .S0(ad[4])
);
MUX2 mux_inst_120 (
  .O(dout[120]),
  .I0(ram16s_inst_30_dout[120]),
  .I1(ram16s_inst_94_dout[120]),
  .S0(ad[4])
);
MUX2 mux_inst_121 (
  .O(dout[121]),
  .I0(ram16s_inst_30_dout[121]),
  .I1(ram16s_inst_94_dout[121]),
  .S0(ad[4])
);
MUX2 mux_inst_122 (
  .O(dout[122]),
  .I0(ram16s_inst_30_dout[122]),
  .I1(ram16s_inst_94_dout[122]),
  .S0(ad[4])
);
MUX2 mux_inst_123 (
  .O(dout[123]),
  .I0(ram16s_inst_30_dout[123]),
  .I1(ram16s_inst_94_dout[123]),
  .S0(ad[4])
);
MUX2 mux_inst_124 (
  .O(dout[124]),
  .I0(ram16s_inst_31_dout[124]),
  .I1(ram16s_inst_95_dout[124]),
  .S0(ad[4])
);
MUX2 mux_inst_125 (
  .O(dout[125]),
  .I0(ram16s_inst_31_dout[125]),
  .I1(ram16s_inst_95_dout[125]),
  .S0(ad[4])
);
MUX2 mux_inst_126 (
  .O(dout[126]),
  .I0(ram16s_inst_31_dout[126]),
  .I1(ram16s_inst_95_dout[126]),
  .S0(ad[4])
);
MUX2 mux_inst_127 (
  .O(dout[127]),
  .I0(ram16s_inst_31_dout[127]),
  .I1(ram16s_inst_95_dout[127]),
  .S0(ad[4])
);
MUX2 mux_inst_128 (
  .O(dout[128]),
  .I0(ram16s_inst_32_dout[128]),
  .I1(ram16s_inst_96_dout[128]),
  .S0(ad[4])
);
MUX2 mux_inst_129 (
  .O(dout[129]),
  .I0(ram16s_inst_32_dout[129]),
  .I1(ram16s_inst_96_dout[129]),
  .S0(ad[4])
);
MUX2 mux_inst_130 (
  .O(dout[130]),
  .I0(ram16s_inst_32_dout[130]),
  .I1(ram16s_inst_96_dout[130]),
  .S0(ad[4])
);
MUX2 mux_inst_131 (
  .O(dout[131]),
  .I0(ram16s_inst_32_dout[131]),
  .I1(ram16s_inst_96_dout[131]),
  .S0(ad[4])
);
MUX2 mux_inst_132 (
  .O(dout[132]),
  .I0(ram16s_inst_33_dout[132]),
  .I1(ram16s_inst_97_dout[132]),
  .S0(ad[4])
);
MUX2 mux_inst_133 (
  .O(dout[133]),
  .I0(ram16s_inst_33_dout[133]),
  .I1(ram16s_inst_97_dout[133]),
  .S0(ad[4])
);
MUX2 mux_inst_134 (
  .O(dout[134]),
  .I0(ram16s_inst_33_dout[134]),
  .I1(ram16s_inst_97_dout[134]),
  .S0(ad[4])
);
MUX2 mux_inst_135 (
  .O(dout[135]),
  .I0(ram16s_inst_33_dout[135]),
  .I1(ram16s_inst_97_dout[135]),
  .S0(ad[4])
);
MUX2 mux_inst_136 (
  .O(dout[136]),
  .I0(ram16s_inst_34_dout[136]),
  .I1(ram16s_inst_98_dout[136]),
  .S0(ad[4])
);
MUX2 mux_inst_137 (
  .O(dout[137]),
  .I0(ram16s_inst_34_dout[137]),
  .I1(ram16s_inst_98_dout[137]),
  .S0(ad[4])
);
MUX2 mux_inst_138 (
  .O(dout[138]),
  .I0(ram16s_inst_34_dout[138]),
  .I1(ram16s_inst_98_dout[138]),
  .S0(ad[4])
);
MUX2 mux_inst_139 (
  .O(dout[139]),
  .I0(ram16s_inst_34_dout[139]),
  .I1(ram16s_inst_98_dout[139]),
  .S0(ad[4])
);
MUX2 mux_inst_140 (
  .O(dout[140]),
  .I0(ram16s_inst_35_dout[140]),
  .I1(ram16s_inst_99_dout[140]),
  .S0(ad[4])
);
MUX2 mux_inst_141 (
  .O(dout[141]),
  .I0(ram16s_inst_35_dout[141]),
  .I1(ram16s_inst_99_dout[141]),
  .S0(ad[4])
);
MUX2 mux_inst_142 (
  .O(dout[142]),
  .I0(ram16s_inst_35_dout[142]),
  .I1(ram16s_inst_99_dout[142]),
  .S0(ad[4])
);
MUX2 mux_inst_143 (
  .O(dout[143]),
  .I0(ram16s_inst_35_dout[143]),
  .I1(ram16s_inst_99_dout[143]),
  .S0(ad[4])
);
MUX2 mux_inst_144 (
  .O(dout[144]),
  .I0(ram16s_inst_36_dout[144]),
  .I1(ram16s_inst_100_dout[144]),
  .S0(ad[4])
);
MUX2 mux_inst_145 (
  .O(dout[145]),
  .I0(ram16s_inst_36_dout[145]),
  .I1(ram16s_inst_100_dout[145]),
  .S0(ad[4])
);
MUX2 mux_inst_146 (
  .O(dout[146]),
  .I0(ram16s_inst_36_dout[146]),
  .I1(ram16s_inst_100_dout[146]),
  .S0(ad[4])
);
MUX2 mux_inst_147 (
  .O(dout[147]),
  .I0(ram16s_inst_36_dout[147]),
  .I1(ram16s_inst_100_dout[147]),
  .S0(ad[4])
);
MUX2 mux_inst_148 (
  .O(dout[148]),
  .I0(ram16s_inst_37_dout[148]),
  .I1(ram16s_inst_101_dout[148]),
  .S0(ad[4])
);
MUX2 mux_inst_149 (
  .O(dout[149]),
  .I0(ram16s_inst_37_dout[149]),
  .I1(ram16s_inst_101_dout[149]),
  .S0(ad[4])
);
MUX2 mux_inst_150 (
  .O(dout[150]),
  .I0(ram16s_inst_37_dout[150]),
  .I1(ram16s_inst_101_dout[150]),
  .S0(ad[4])
);
MUX2 mux_inst_151 (
  .O(dout[151]),
  .I0(ram16s_inst_37_dout[151]),
  .I1(ram16s_inst_101_dout[151]),
  .S0(ad[4])
);
MUX2 mux_inst_152 (
  .O(dout[152]),
  .I0(ram16s_inst_38_dout[152]),
  .I1(ram16s_inst_102_dout[152]),
  .S0(ad[4])
);
MUX2 mux_inst_153 (
  .O(dout[153]),
  .I0(ram16s_inst_38_dout[153]),
  .I1(ram16s_inst_102_dout[153]),
  .S0(ad[4])
);
MUX2 mux_inst_154 (
  .O(dout[154]),
  .I0(ram16s_inst_38_dout[154]),
  .I1(ram16s_inst_102_dout[154]),
  .S0(ad[4])
);
MUX2 mux_inst_155 (
  .O(dout[155]),
  .I0(ram16s_inst_38_dout[155]),
  .I1(ram16s_inst_102_dout[155]),
  .S0(ad[4])
);
MUX2 mux_inst_156 (
  .O(dout[156]),
  .I0(ram16s_inst_39_dout[156]),
  .I1(ram16s_inst_103_dout[156]),
  .S0(ad[4])
);
MUX2 mux_inst_157 (
  .O(dout[157]),
  .I0(ram16s_inst_39_dout[157]),
  .I1(ram16s_inst_103_dout[157]),
  .S0(ad[4])
);
MUX2 mux_inst_158 (
  .O(dout[158]),
  .I0(ram16s_inst_39_dout[158]),
  .I1(ram16s_inst_103_dout[158]),
  .S0(ad[4])
);
MUX2 mux_inst_159 (
  .O(dout[159]),
  .I0(ram16s_inst_39_dout[159]),
  .I1(ram16s_inst_103_dout[159]),
  .S0(ad[4])
);
MUX2 mux_inst_160 (
  .O(dout[160]),
  .I0(ram16s_inst_40_dout[160]),
  .I1(ram16s_inst_104_dout[160]),
  .S0(ad[4])
);
MUX2 mux_inst_161 (
  .O(dout[161]),
  .I0(ram16s_inst_40_dout[161]),
  .I1(ram16s_inst_104_dout[161]),
  .S0(ad[4])
);
MUX2 mux_inst_162 (
  .O(dout[162]),
  .I0(ram16s_inst_40_dout[162]),
  .I1(ram16s_inst_104_dout[162]),
  .S0(ad[4])
);
MUX2 mux_inst_163 (
  .O(dout[163]),
  .I0(ram16s_inst_40_dout[163]),
  .I1(ram16s_inst_104_dout[163]),
  .S0(ad[4])
);
MUX2 mux_inst_164 (
  .O(dout[164]),
  .I0(ram16s_inst_41_dout[164]),
  .I1(ram16s_inst_105_dout[164]),
  .S0(ad[4])
);
MUX2 mux_inst_165 (
  .O(dout[165]),
  .I0(ram16s_inst_41_dout[165]),
  .I1(ram16s_inst_105_dout[165]),
  .S0(ad[4])
);
MUX2 mux_inst_166 (
  .O(dout[166]),
  .I0(ram16s_inst_41_dout[166]),
  .I1(ram16s_inst_105_dout[166]),
  .S0(ad[4])
);
MUX2 mux_inst_167 (
  .O(dout[167]),
  .I0(ram16s_inst_41_dout[167]),
  .I1(ram16s_inst_105_dout[167]),
  .S0(ad[4])
);
MUX2 mux_inst_168 (
  .O(dout[168]),
  .I0(ram16s_inst_42_dout[168]),
  .I1(ram16s_inst_106_dout[168]),
  .S0(ad[4])
);
MUX2 mux_inst_169 (
  .O(dout[169]),
  .I0(ram16s_inst_42_dout[169]),
  .I1(ram16s_inst_106_dout[169]),
  .S0(ad[4])
);
MUX2 mux_inst_170 (
  .O(dout[170]),
  .I0(ram16s_inst_42_dout[170]),
  .I1(ram16s_inst_106_dout[170]),
  .S0(ad[4])
);
MUX2 mux_inst_171 (
  .O(dout[171]),
  .I0(ram16s_inst_42_dout[171]),
  .I1(ram16s_inst_106_dout[171]),
  .S0(ad[4])
);
MUX2 mux_inst_172 (
  .O(dout[172]),
  .I0(ram16s_inst_43_dout[172]),
  .I1(ram16s_inst_107_dout[172]),
  .S0(ad[4])
);
MUX2 mux_inst_173 (
  .O(dout[173]),
  .I0(ram16s_inst_43_dout[173]),
  .I1(ram16s_inst_107_dout[173]),
  .S0(ad[4])
);
MUX2 mux_inst_174 (
  .O(dout[174]),
  .I0(ram16s_inst_43_dout[174]),
  .I1(ram16s_inst_107_dout[174]),
  .S0(ad[4])
);
MUX2 mux_inst_175 (
  .O(dout[175]),
  .I0(ram16s_inst_43_dout[175]),
  .I1(ram16s_inst_107_dout[175]),
  .S0(ad[4])
);
MUX2 mux_inst_176 (
  .O(dout[176]),
  .I0(ram16s_inst_44_dout[176]),
  .I1(ram16s_inst_108_dout[176]),
  .S0(ad[4])
);
MUX2 mux_inst_177 (
  .O(dout[177]),
  .I0(ram16s_inst_44_dout[177]),
  .I1(ram16s_inst_108_dout[177]),
  .S0(ad[4])
);
MUX2 mux_inst_178 (
  .O(dout[178]),
  .I0(ram16s_inst_44_dout[178]),
  .I1(ram16s_inst_108_dout[178]),
  .S0(ad[4])
);
MUX2 mux_inst_179 (
  .O(dout[179]),
  .I0(ram16s_inst_44_dout[179]),
  .I1(ram16s_inst_108_dout[179]),
  .S0(ad[4])
);
MUX2 mux_inst_180 (
  .O(dout[180]),
  .I0(ram16s_inst_45_dout[180]),
  .I1(ram16s_inst_109_dout[180]),
  .S0(ad[4])
);
MUX2 mux_inst_181 (
  .O(dout[181]),
  .I0(ram16s_inst_45_dout[181]),
  .I1(ram16s_inst_109_dout[181]),
  .S0(ad[4])
);
MUX2 mux_inst_182 (
  .O(dout[182]),
  .I0(ram16s_inst_45_dout[182]),
  .I1(ram16s_inst_109_dout[182]),
  .S0(ad[4])
);
MUX2 mux_inst_183 (
  .O(dout[183]),
  .I0(ram16s_inst_45_dout[183]),
  .I1(ram16s_inst_109_dout[183]),
  .S0(ad[4])
);
MUX2 mux_inst_184 (
  .O(dout[184]),
  .I0(ram16s_inst_46_dout[184]),
  .I1(ram16s_inst_110_dout[184]),
  .S0(ad[4])
);
MUX2 mux_inst_185 (
  .O(dout[185]),
  .I0(ram16s_inst_46_dout[185]),
  .I1(ram16s_inst_110_dout[185]),
  .S0(ad[4])
);
MUX2 mux_inst_186 (
  .O(dout[186]),
  .I0(ram16s_inst_46_dout[186]),
  .I1(ram16s_inst_110_dout[186]),
  .S0(ad[4])
);
MUX2 mux_inst_187 (
  .O(dout[187]),
  .I0(ram16s_inst_46_dout[187]),
  .I1(ram16s_inst_110_dout[187]),
  .S0(ad[4])
);
MUX2 mux_inst_188 (
  .O(dout[188]),
  .I0(ram16s_inst_47_dout[188]),
  .I1(ram16s_inst_111_dout[188]),
  .S0(ad[4])
);
MUX2 mux_inst_189 (
  .O(dout[189]),
  .I0(ram16s_inst_47_dout[189]),
  .I1(ram16s_inst_111_dout[189]),
  .S0(ad[4])
);
MUX2 mux_inst_190 (
  .O(dout[190]),
  .I0(ram16s_inst_47_dout[190]),
  .I1(ram16s_inst_111_dout[190]),
  .S0(ad[4])
);
MUX2 mux_inst_191 (
  .O(dout[191]),
  .I0(ram16s_inst_47_dout[191]),
  .I1(ram16s_inst_111_dout[191]),
  .S0(ad[4])
);
MUX2 mux_inst_192 (
  .O(dout[192]),
  .I0(ram16s_inst_48_dout[192]),
  .I1(ram16s_inst_112_dout[192]),
  .S0(ad[4])
);
MUX2 mux_inst_193 (
  .O(dout[193]),
  .I0(ram16s_inst_48_dout[193]),
  .I1(ram16s_inst_112_dout[193]),
  .S0(ad[4])
);
MUX2 mux_inst_194 (
  .O(dout[194]),
  .I0(ram16s_inst_48_dout[194]),
  .I1(ram16s_inst_112_dout[194]),
  .S0(ad[4])
);
MUX2 mux_inst_195 (
  .O(dout[195]),
  .I0(ram16s_inst_48_dout[195]),
  .I1(ram16s_inst_112_dout[195]),
  .S0(ad[4])
);
MUX2 mux_inst_196 (
  .O(dout[196]),
  .I0(ram16s_inst_49_dout[196]),
  .I1(ram16s_inst_113_dout[196]),
  .S0(ad[4])
);
MUX2 mux_inst_197 (
  .O(dout[197]),
  .I0(ram16s_inst_49_dout[197]),
  .I1(ram16s_inst_113_dout[197]),
  .S0(ad[4])
);
MUX2 mux_inst_198 (
  .O(dout[198]),
  .I0(ram16s_inst_49_dout[198]),
  .I1(ram16s_inst_113_dout[198]),
  .S0(ad[4])
);
MUX2 mux_inst_199 (
  .O(dout[199]),
  .I0(ram16s_inst_49_dout[199]),
  .I1(ram16s_inst_113_dout[199]),
  .S0(ad[4])
);
MUX2 mux_inst_200 (
  .O(dout[200]),
  .I0(ram16s_inst_50_dout[200]),
  .I1(ram16s_inst_114_dout[200]),
  .S0(ad[4])
);
MUX2 mux_inst_201 (
  .O(dout[201]),
  .I0(ram16s_inst_50_dout[201]),
  .I1(ram16s_inst_114_dout[201]),
  .S0(ad[4])
);
MUX2 mux_inst_202 (
  .O(dout[202]),
  .I0(ram16s_inst_50_dout[202]),
  .I1(ram16s_inst_114_dout[202]),
  .S0(ad[4])
);
MUX2 mux_inst_203 (
  .O(dout[203]),
  .I0(ram16s_inst_50_dout[203]),
  .I1(ram16s_inst_114_dout[203]),
  .S0(ad[4])
);
MUX2 mux_inst_204 (
  .O(dout[204]),
  .I0(ram16s_inst_51_dout[204]),
  .I1(ram16s_inst_115_dout[204]),
  .S0(ad[4])
);
MUX2 mux_inst_205 (
  .O(dout[205]),
  .I0(ram16s_inst_51_dout[205]),
  .I1(ram16s_inst_115_dout[205]),
  .S0(ad[4])
);
MUX2 mux_inst_206 (
  .O(dout[206]),
  .I0(ram16s_inst_51_dout[206]),
  .I1(ram16s_inst_115_dout[206]),
  .S0(ad[4])
);
MUX2 mux_inst_207 (
  .O(dout[207]),
  .I0(ram16s_inst_51_dout[207]),
  .I1(ram16s_inst_115_dout[207]),
  .S0(ad[4])
);
MUX2 mux_inst_208 (
  .O(dout[208]),
  .I0(ram16s_inst_52_dout[208]),
  .I1(ram16s_inst_116_dout[208]),
  .S0(ad[4])
);
MUX2 mux_inst_209 (
  .O(dout[209]),
  .I0(ram16s_inst_52_dout[209]),
  .I1(ram16s_inst_116_dout[209]),
  .S0(ad[4])
);
MUX2 mux_inst_210 (
  .O(dout[210]),
  .I0(ram16s_inst_52_dout[210]),
  .I1(ram16s_inst_116_dout[210]),
  .S0(ad[4])
);
MUX2 mux_inst_211 (
  .O(dout[211]),
  .I0(ram16s_inst_52_dout[211]),
  .I1(ram16s_inst_116_dout[211]),
  .S0(ad[4])
);
MUX2 mux_inst_212 (
  .O(dout[212]),
  .I0(ram16s_inst_53_dout[212]),
  .I1(ram16s_inst_117_dout[212]),
  .S0(ad[4])
);
MUX2 mux_inst_213 (
  .O(dout[213]),
  .I0(ram16s_inst_53_dout[213]),
  .I1(ram16s_inst_117_dout[213]),
  .S0(ad[4])
);
MUX2 mux_inst_214 (
  .O(dout[214]),
  .I0(ram16s_inst_53_dout[214]),
  .I1(ram16s_inst_117_dout[214]),
  .S0(ad[4])
);
MUX2 mux_inst_215 (
  .O(dout[215]),
  .I0(ram16s_inst_53_dout[215]),
  .I1(ram16s_inst_117_dout[215]),
  .S0(ad[4])
);
MUX2 mux_inst_216 (
  .O(dout[216]),
  .I0(ram16s_inst_54_dout[216]),
  .I1(ram16s_inst_118_dout[216]),
  .S0(ad[4])
);
MUX2 mux_inst_217 (
  .O(dout[217]),
  .I0(ram16s_inst_54_dout[217]),
  .I1(ram16s_inst_118_dout[217]),
  .S0(ad[4])
);
MUX2 mux_inst_218 (
  .O(dout[218]),
  .I0(ram16s_inst_54_dout[218]),
  .I1(ram16s_inst_118_dout[218]),
  .S0(ad[4])
);
MUX2 mux_inst_219 (
  .O(dout[219]),
  .I0(ram16s_inst_54_dout[219]),
  .I1(ram16s_inst_118_dout[219]),
  .S0(ad[4])
);
MUX2 mux_inst_220 (
  .O(dout[220]),
  .I0(ram16s_inst_55_dout[220]),
  .I1(ram16s_inst_119_dout[220]),
  .S0(ad[4])
);
MUX2 mux_inst_221 (
  .O(dout[221]),
  .I0(ram16s_inst_55_dout[221]),
  .I1(ram16s_inst_119_dout[221]),
  .S0(ad[4])
);
MUX2 mux_inst_222 (
  .O(dout[222]),
  .I0(ram16s_inst_55_dout[222]),
  .I1(ram16s_inst_119_dout[222]),
  .S0(ad[4])
);
MUX2 mux_inst_223 (
  .O(dout[223]),
  .I0(ram16s_inst_55_dout[223]),
  .I1(ram16s_inst_119_dout[223]),
  .S0(ad[4])
);
MUX2 mux_inst_224 (
  .O(dout[224]),
  .I0(ram16s_inst_56_dout[224]),
  .I1(ram16s_inst_120_dout[224]),
  .S0(ad[4])
);
MUX2 mux_inst_225 (
  .O(dout[225]),
  .I0(ram16s_inst_56_dout[225]),
  .I1(ram16s_inst_120_dout[225]),
  .S0(ad[4])
);
MUX2 mux_inst_226 (
  .O(dout[226]),
  .I0(ram16s_inst_56_dout[226]),
  .I1(ram16s_inst_120_dout[226]),
  .S0(ad[4])
);
MUX2 mux_inst_227 (
  .O(dout[227]),
  .I0(ram16s_inst_56_dout[227]),
  .I1(ram16s_inst_120_dout[227]),
  .S0(ad[4])
);
MUX2 mux_inst_228 (
  .O(dout[228]),
  .I0(ram16s_inst_57_dout[228]),
  .I1(ram16s_inst_121_dout[228]),
  .S0(ad[4])
);
MUX2 mux_inst_229 (
  .O(dout[229]),
  .I0(ram16s_inst_57_dout[229]),
  .I1(ram16s_inst_121_dout[229]),
  .S0(ad[4])
);
MUX2 mux_inst_230 (
  .O(dout[230]),
  .I0(ram16s_inst_57_dout[230]),
  .I1(ram16s_inst_121_dout[230]),
  .S0(ad[4])
);
MUX2 mux_inst_231 (
  .O(dout[231]),
  .I0(ram16s_inst_57_dout[231]),
  .I1(ram16s_inst_121_dout[231]),
  .S0(ad[4])
);
MUX2 mux_inst_232 (
  .O(dout[232]),
  .I0(ram16s_inst_58_dout[232]),
  .I1(ram16s_inst_122_dout[232]),
  .S0(ad[4])
);
MUX2 mux_inst_233 (
  .O(dout[233]),
  .I0(ram16s_inst_58_dout[233]),
  .I1(ram16s_inst_122_dout[233]),
  .S0(ad[4])
);
MUX2 mux_inst_234 (
  .O(dout[234]),
  .I0(ram16s_inst_58_dout[234]),
  .I1(ram16s_inst_122_dout[234]),
  .S0(ad[4])
);
MUX2 mux_inst_235 (
  .O(dout[235]),
  .I0(ram16s_inst_58_dout[235]),
  .I1(ram16s_inst_122_dout[235]),
  .S0(ad[4])
);
MUX2 mux_inst_236 (
  .O(dout[236]),
  .I0(ram16s_inst_59_dout[236]),
  .I1(ram16s_inst_123_dout[236]),
  .S0(ad[4])
);
MUX2 mux_inst_237 (
  .O(dout[237]),
  .I0(ram16s_inst_59_dout[237]),
  .I1(ram16s_inst_123_dout[237]),
  .S0(ad[4])
);
MUX2 mux_inst_238 (
  .O(dout[238]),
  .I0(ram16s_inst_59_dout[238]),
  .I1(ram16s_inst_123_dout[238]),
  .S0(ad[4])
);
MUX2 mux_inst_239 (
  .O(dout[239]),
  .I0(ram16s_inst_59_dout[239]),
  .I1(ram16s_inst_123_dout[239]),
  .S0(ad[4])
);
MUX2 mux_inst_240 (
  .O(dout[240]),
  .I0(ram16s_inst_60_dout[240]),
  .I1(ram16s_inst_124_dout[240]),
  .S0(ad[4])
);
MUX2 mux_inst_241 (
  .O(dout[241]),
  .I0(ram16s_inst_60_dout[241]),
  .I1(ram16s_inst_124_dout[241]),
  .S0(ad[4])
);
MUX2 mux_inst_242 (
  .O(dout[242]),
  .I0(ram16s_inst_60_dout[242]),
  .I1(ram16s_inst_124_dout[242]),
  .S0(ad[4])
);
MUX2 mux_inst_243 (
  .O(dout[243]),
  .I0(ram16s_inst_60_dout[243]),
  .I1(ram16s_inst_124_dout[243]),
  .S0(ad[4])
);
MUX2 mux_inst_244 (
  .O(dout[244]),
  .I0(ram16s_inst_61_dout[244]),
  .I1(ram16s_inst_125_dout[244]),
  .S0(ad[4])
);
MUX2 mux_inst_245 (
  .O(dout[245]),
  .I0(ram16s_inst_61_dout[245]),
  .I1(ram16s_inst_125_dout[245]),
  .S0(ad[4])
);
MUX2 mux_inst_246 (
  .O(dout[246]),
  .I0(ram16s_inst_61_dout[246]),
  .I1(ram16s_inst_125_dout[246]),
  .S0(ad[4])
);
MUX2 mux_inst_247 (
  .O(dout[247]),
  .I0(ram16s_inst_61_dout[247]),
  .I1(ram16s_inst_125_dout[247]),
  .S0(ad[4])
);
MUX2 mux_inst_248 (
  .O(dout[248]),
  .I0(ram16s_inst_62_dout[248]),
  .I1(ram16s_inst_126_dout[248]),
  .S0(ad[4])
);
MUX2 mux_inst_249 (
  .O(dout[249]),
  .I0(ram16s_inst_62_dout[249]),
  .I1(ram16s_inst_126_dout[249]),
  .S0(ad[4])
);
MUX2 mux_inst_250 (
  .O(dout[250]),
  .I0(ram16s_inst_62_dout[250]),
  .I1(ram16s_inst_126_dout[250]),
  .S0(ad[4])
);
MUX2 mux_inst_251 (
  .O(dout[251]),
  .I0(ram16s_inst_62_dout[251]),
  .I1(ram16s_inst_126_dout[251]),
  .S0(ad[4])
);
MUX2 mux_inst_252 (
  .O(dout[252]),
  .I0(ram16s_inst_63_dout[252]),
  .I1(ram16s_inst_127_dout[252]),
  .S0(ad[4])
);
MUX2 mux_inst_253 (
  .O(dout[253]),
  .I0(ram16s_inst_63_dout[253]),
  .I1(ram16s_inst_127_dout[253]),
  .S0(ad[4])
);
MUX2 mux_inst_254 (
  .O(dout[254]),
  .I0(ram16s_inst_63_dout[254]),
  .I1(ram16s_inst_127_dout[254]),
  .S0(ad[4])
);
MUX2 mux_inst_255 (
  .O(dout[255]),
  .I0(ram16s_inst_63_dout[255]),
  .I1(ram16s_inst_127_dout[255]),
  .S0(ad[4])
);
endmodule //Gowin_RAM16S
