// Instantiation of core and cache memory
