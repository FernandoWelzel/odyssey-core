// Processor core
module core #(
    parameter DATA_WIDTH = 32
)
(
    input  logic clk,
    input  logic rst
);

// Fetch instantiation
// Decode instantiation
// ALU instantiation
// Register file instantiation
// LSU instantiation

endmodule
