// Processor load and store unit
module lsu #(
    parameter DATA_WIDTH = 32
)
(
    input  logic clk,
    input  logic rst
);

endmodule
