// Processor decode unit
module decode #(
    parameter DATA_WIDTH = 32
)
(
    input  logic clk,
    input  logic rst
);

endmodule
