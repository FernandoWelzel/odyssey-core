// Processor register file
module register_file #(
    parameter REGISTERS = 32
)
(
    input  logic clk,
    input  logic rst
);

endmodule
